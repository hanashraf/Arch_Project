library verilog;
use verilog.vl_types.all;
entity testbench_tx is
end testbench_tx;
