library verilog;
use verilog.vl_types.all;
entity testbench_bd is
end testbench_bd;
