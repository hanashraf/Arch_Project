library verilog;
use verilog.vl_types.all;
entity testbench_slave is
end testbench_slave;
