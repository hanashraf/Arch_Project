library verilog;
use verilog.vl_types.all;
entity testbench_rx is
end testbench_rx;
