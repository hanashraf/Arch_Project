library verilog;
use verilog.vl_types.all;
entity testbench_oversampling is
end testbench_oversampling;
