module testbench_rx();
  // Declare input and output signals for the MUT
  reg clk;
  reg rst;
  reg rxd;
  wire [7:0] rec_data_out;
  wire rec_valid_out;

  // Instantiate the MUT
  rx MUT (
    .clk(clk),
    .rst(rst),
    .rxd(rxd),
    .rec_data_out(rec_data_out),
    .rec_valid_out(rec_valid_out)
  );

  // Initialize input signals and registers
  initial begin
    clk = 0;
    rst = 1;
    rxd = 0;
    #10 rst = 0;
  end

  // Apply stimuli to the MUT and observe the output responses
  always begin
    #5 clk = ~clk;
  end

  // Print out input and output signals
  initial begin
    $monitor("rxd=%d rec_data=%d rec_valid=%d", rxd, rec_data_out, rec_valid_out);
  end

   // Test case: receive multiple data words
  initial begin
    rxd = 1;
    #100; rxd = 0;
    #40; rxd = 1;
    #40; rxd = 0;
    #40; rxd = 1;
    #40; rxd = 0;
  end

endmodule



